--##########################################################################################--
--########### GŁÓWNI AUTORZY KODU DO IMPEMENTACJI: JAKUB OBACZ, MICHAL POPEK ###############--
--############## AUTORZY TESTÓW: MATEUSZ WOLAK, WIKTOR BAJEWSKI, JAKUB OBACZ ###############--
--##########################################################################################--
library IEEE;
use IEEE.STD_LOGIC_1164.all;

package whitelion is

        type regdatatype is array(15 downto 0) of std_logic_vector(7 downto 0);
        type regwritetype is array(15 downto 0) of std_logic;

end whitelion;

package body whitelion is
end whitelion;
